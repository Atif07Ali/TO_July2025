* Equivalent circuit model for E:\touchstone_files\42p.ckt
.SUBCKT 42p po1 po2
Vsp1 po1 p1 0
Vsr1 p1 pr1 0
Rp1 pr1 0 50
Ru1 u1 0 50
Fr1 u1 0 Vsr1 -1
Fu1 u1 0 Vsp1 -1
Ry1 y1 0 1
Gy1 p1 0 y1 0 -0.02
Vsp2 po2 p2 0
Vsr2 p2 pr2 0
Rp2 pr2 0 50
Ru2 u2 0 50
Fr2 u2 0 Vsr2 -1
Fu2 u2 0 Vsp2 -1
Ry2 y2 0 1
Gy2 p2 0 y2 0 -0.02
Rx1 x1 0 1
Fxc1_2 x1 0 Vx2 0.0506033419001637
Cx1 x1 xm1 3.42335591038431e-13
Vx1 xm1 0 0
Gx1_1 x1 0 u1 0 -0.0837230038088886
Rx2 x2 0 1
Fxc2_1 x2 0 Vx1 -9.08119096919164
Cx2 x2 xm2 3.42335591038431e-13
Vx2 xm2 0 0
Gx2_1 x2 0 u1 0 0.760304586102876
Rx3 x3 0 1
Fxc3_4 x3 0 Vx4 3.36907918673722
Cx3 x3 xm3 1.14997202900161e-13
Vx3 xm3 0 0
Gx3_1 x3 0 u1 0 -0.171097604429355
Rx4 x4 0 1
Fxc4_3 x4 0 Vx3 -1.85350835822414
Cx4 x4 xm4 1.14997202900161e-13
Vx4 xm4 0 0
Gx4_1 x4 0 u1 0 0.317130839881936
Rx5 x5 0 1
Cx5 x5 0 6.34424328985755e-12
Gx5_1 x5 0 u1 0 -0.00761686241004208
Rx6 x6 0 1
Fxc6_7 x6 0 Vx7 0.0505300699899194
Cx6 x6 xm6 3.42335591038431e-13
Vx6 xm6 0 0
Gx6_2 x6 0 u2 0 -0.0836063384059733
Rx7 x7 0 1
Fxc7_6 x7 0 Vx6 -9.09435929074232
Cx7 x7 xm7 3.42335591038431e-13
Vx7 xm7 0 0
Gx7_2 x7 0 u2 0 0.760346080447309
Rx8 x8 0 1
Fxc8_9 x8 0 Vx9 3.36807785871027
Cx8 x8 xm8 1.14997202900161e-13
Vx8 xm8 0 0
Gx8_2 x8 0 u2 0 -0.171071010729707
Rx9 x9 0 1
Fxc9_8 x9 0 Vx8 -1.85405940542231
Cx9 x9 xm9 1.14997202900161e-13
Vx9 xm9 0 0
Gx9_2 x9 0 u2 0 0.317175816438514
Rx10 x10 0 1
Cx10 x10 0 6.34424328985755e-12
Gx10_2 x10 0 u2 0 -0.00762042787610135
Gyc1_1 y1 0 x1 0 0.660729716006035
Gyc1_2 y1 0 x2 0 0.0831777594333287
Gyc1_3 y1 0 x3 0 -0.051735576347353
Gyc1_4 y1 0 x4 0 -0.0320154148016977
Gyc1_5 y1 0 x5 0 0.478815278418924
Gyc1_6 y1 0 x6 0 -1
Gyc1_7 y1 0 x7 0 1
Gyc1_8 y1 0 x8 0 1
Gyc1_9 y1 0 x9 0 1
Gyc1_10 y1 0 x10 0 -1
Gyc2_1 y2 0 x1 0 -1
Gyc2_2 y2 0 x2 0 1
Gyc2_3 y2 0 x3 0 1
Gyc2_4 y2 0 x4 0 1
Gyc2_5 y2 0 x5 0 -1
Gyc2_6 y2 0 x6 0 0.634392213787007
Gyc2_7 y2 0 x7 0 0.082279060093136
Gyc2_8 y2 0 x8 0 -0.0512941134164529
Gyc2_9 y2 0 x9 0 -0.0369413839527659
Gyc2_10 y2 0 x10 0 0.473691375648657
.ENDS
