* Equivalent circuit model for E:\touchstone_files\choke_first1.ckt
.SUBCKT choke_first1 po1 po2
Vsp1 po1 p1 0
Vsr1 p1 pr1 0
Rp1 pr1 0 50
Ru1 u1 0 50
Fr1 u1 0 Vsr1 -1
Fu1 u1 0 Vsp1 -1
Ry1 y1 0 1
Gy1 p1 0 y1 0 -0.02
Vsp2 po2 p2 0
Vsr2 p2 pr2 0
Rp2 pr2 0 50
Ru2 u2 0 50
Fr2 u2 0 Vsr2 -1
Fu2 u2 0 Vsp2 -1
Ry2 y2 0 1
Gy2 p2 0 y2 0 -0.02
Rx1 x1 0 1
Fxc1_2 x1 0 Vx2 0.101995236600397
Cx1 x1 xm1 3.69242380877071e-13
Vx1 xm1 0 0
Gx1_1 x1 0 u1 0 -2.33209763814394
Rx2 x2 0 1
Fxc2_1 x2 0 Vx1 -3.61108727128201
Cx2 x2 xm2 3.69242380877071e-13
Vx2 xm2 0 0
Gx2_1 x2 0 u1 0 8.42140809648841
Rx3 x3 0 1
Fxc3_4 x3 0 Vx4 5.29536141445428
Cx3 x3 xm3 1.07756536529339e-13
Vx3 xm3 0 0
Gx3_1 x3 0 u1 0 -1.04743590328075
Rx4 x4 0 1
Fxc4_3 x4 0 Vx3 -1.02776588658002
Cx4 x4 xm4 1.07756536529339e-13
Vx4 xm4 0 0
Gx4_1 x4 0 u1 0 1.07651888977109
Rx5 x5 0 1
Fxc5_6 x5 0 Vx6 0.428667781676471
Cx5 x5 xm5 1.10864231314785e-12
Vx5 xm5 0 0
Gx5_1 x5 0 u1 0 -4.40084921808134
Rx6 x6 0 1
Fxc6_5 x6 0 Vx5 -0.441808922439799
Cx6 x6 xm6 1.10864231314785e-12
Vx6 xm6 0 0
Gx6_1 x6 0 u1 0 1.94433445086055
Rx7 x7 0 1
Fxc7_8 x7 0 Vx8 1.63850227458527
Cx7 x7 xm7 3.10221523673382e-13
Vx7 xm7 0 0
Gx7_1 x7 0 u1 0 -0.202614926478493
Rx8 x8 0 1
Fxc8_7 x8 0 Vx7 -2.27068857006175
Cx8 x8 xm8 3.10221523673382e-13
Vx8 xm8 0 0
Gx8_1 x8 0 u1 0 0.460075397678615
Rx9 x9 0 1
Fxc9_10 x9 0 Vx10 4.82487580664991
Cx9 x9 xm9 8.39178096976935e-14
Vx9 xm9 0 0
Gx9_1 x9 0 u1 0 -0.0103038151219182
Rx10 x10 0 1
Fxc10_9 x10 0 Vx9 -7.17961729578961
Cx10 x10 xm10 8.39178096976935e-14
Vx10 xm10 0 0
Gx10_1 x10 0 u1 0 0.0739774492619424
Rx11 x11 0 1
Cx11 x11 0 3.05463655648388e-12
Gx11_1 x11 0 u1 0 -2.83630053852568
Rx12 x12 0 1
Fxc12_13 x12 0 Vx13 0.201636688353947
Cx12 x12 xm12 3.69242380877071e-13
Vx12 xm12 0 0
Gx12_2 x12 0 u2 0 -2.61120485734652
Rx13 x13 0 1
Fxc13_12 x13 0 Vx12 -1.82662046091813
Cx13 x13 xm13 3.69242380877071e-13
Vx13 xm13 0 0
Gx13_2 x13 0 u2 0 4.76968022007795
Rx14 x14 0 1
Fxc14_15 x14 0 Vx15 1.44819583555059
Cx14 x14 xm14 1.07756536529339e-13
Vx14 xm14 0 0
Gx14_2 x14 0 u2 0 -0.354376395935862
Rx15 x15 0 1
Fxc15_14 x15 0 Vx14 -3.75804962649895
Cx15 x15 xm15 1.07756536529339e-13
Vx15 xm15 0 0
Gx15_2 x15 0 u2 0 1.33176408238681
Rx16 x16 0 1
Fxc16_17 x16 0 Vx17 0.441992282984616
Cx16 x16 xm16 1.10864231314785e-12
Vx16 xm16 0 0
Gx16_2 x16 0 u2 0 -4.31856642795994
Rx17 x17 0 1
Fxc17_16 x17 0 Vx16 -0.428489948802415
Cx17 x17 xm17 1.10864231314785e-12
Vx17 xm17 0 0
Gx17_2 x17 0 u2 0 1.85046230761638
Rx18 x18 0 1
Fxc18_19 x18 0 Vx19 1.58791262650135
Cx18 x18 xm18 3.10221523673382e-13
Vx18 xm18 0 0
Gx18_2 x18 0 u2 0 -0.19170048357859
Rx19 x19 0 1
Fxc19_18 x19 0 Vx18 -2.34303092300386
Cx19 x19 xm19 3.10221523673382e-13
Vx19 xm19 0 0
Gx19_2 x19 0 u2 0 0.44916016097943
Rx20 x20 0 1
Fxc20_21 x20 0 Vx21 4.87371342501607
Cx20 x20 xm20 8.39178096976935e-14
Vx20 xm20 0 0
Gx20_2 x20 0 u2 0 -0.00970566763378732
Rx21 x21 0 1
Fxc21_20 x21 0 Vx20 -7.10767309658677
Cx21 x21 xm21 8.39178096976935e-14
Vx21 xm21 0 0
Gx21_2 x21 0 u2 0 0.0689847127250832
Rx22 x22 0 1
Cx22 x22 0 3.05463655648388e-12
Gx22_2 x22 0 u2 0 -2.74657278375131
Gyc1_1 y1 0 x1 0 -1
Gyc1_2 y1 0 x2 0 -1
Gyc1_3 y1 0 x3 0 1
Gyc1_4 y1 0 x4 0 1
Gyc1_5 y1 0 x5 0 -1
Gyc1_6 y1 0 x6 0 -1
Gyc1_7 y1 0 x7 0 -0.89586625765799
Gyc1_8 y1 0 x8 0 1
Gyc1_9 y1 0 x9 0 0.446025479038402
Gyc1_10 y1 0 x10 0 1
Gyc1_11 y1 0 x11 0 -1
Gyc1_12 y1 0 x12 0 0.129680953382939
Gyc1_13 y1 0 x13 0 -1
Gyc1_14 y1 0 x14 0 1
Gyc1_15 y1 0 x15 0 0.36612337539922
Gyc1_16 y1 0 x16 0 -1
Gyc1_17 y1 0 x17 0 -1
Gyc1_18 y1 0 x18 0 -0.911297558116988
Gyc1_19 y1 0 x19 0 1
Gyc1_20 y1 0 x20 0 0.479147603745794
Gyc1_21 y1 0 x21 0 1
Gyc1_22 y1 0 x22 0 -1
Gyc2_1 y2 0 x1 0 0.759404698095239
Gyc2_2 y2 0 x2 0 -0.0836745333308788
Gyc2_3 y2 0 x3 0 -0.115612005003245
Gyc2_4 y2 0 x4 0 0.200984326811581
Gyc2_5 y2 0 x5 0 -0.420482058449482
Gyc2_6 y2 0 x6 0 -0.750303735134525
Gyc2_7 y2 0 x7 0 -1
Gyc2_8 y2 0 x8 0 -0.142723051145421
Gyc2_9 y2 0 x9 0 -1
Gyc2_10 y2 0 x10 0 0.334006777325338
Gyc2_11 y2 0 x11 0 -0.877832624115024
Gyc2_12 y2 0 x12 0 1
Gyc2_13 y2 0 x13 0 -0.38390462774705
Gyc2_14 y2 0 x14 0 -0.7993745074972
Gyc2_15 y2 0 x15 0 1
Gyc2_16 y2 0 x16 0 -0.379411368345305
Gyc2_17 y2 0 x17 0 -0.74514453520178
Gyc2_18 y2 0 x18 0 -1
Gyc2_19 y2 0 x19 0 -0.133639671598507
Gyc2_20 y2 0 x20 0 -1
Gyc2_21 y2 0 x21 0 0.334951212412435
Gyc2_22 y2 0 x22 0 -0.852650462755582
.ENDS
