* Equivalent circuit model for E:\touchstone_files\outputplane.ckt
.SUBCKT outputplane po1 po2
Vsp1 po1 p1 0
Vsr1 p1 pr1 0
Rp1 pr1 0 50
Ru1 u1 0 50
Fr1 u1 0 Vsr1 -1
Fu1 u1 0 Vsp1 -1
Ry1 y1 0 1
Gy1 p1 0 y1 0 -0.02
Vsp2 po2 p2 0
Vsr2 p2 pr2 0
Rp2 pr2 0 50
Ru2 u2 0 50
Fr2 u2 0 Vsr2 -1
Fu2 u2 0 Vsp2 -1
Ry2 y2 0 1
Gy2 p2 0 y2 0 -0.02
Rx1 x1 0 1
Fxc1_2 x1 0 Vx2 6.77090506944045
Cx1 x1 xm1 1.22121348511033e-13
Vx1 xm1 0 0
Gx1_1 x1 0 u1 0 -0.669904305545353
Rx2 x2 0 1
Fxc2_1 x2 0 Vx1 -0.48231124160245
Cx2 x2 xm2 1.22121348511033e-13
Vx2 xm2 0 0
Gx2_1 x2 0 u1 0 0.323102377362406
Rx3 x3 0 1
Fxc3_4 x3 0 Vx4 0.363120755884473
Cx3 x3 xm3 2.69558380066553e-12
Vx3 xm3 0 0
Gx3_1 x3 0 u1 0 -4.47908785892089
Rx4 x4 0 1
Fxc4_3 x4 0 Vx3 -0.373469152589108
Cx4 x4 xm4 2.69558380066553e-12
Vx4 xm4 0 0
Gx4_1 x4 0 u1 0 1.67280114704335
Rx5 x5 0 1
Fxc5_6 x5 0 Vx6 0.272584774586069
Cx5 x5 xm5 1.3632937533957e-12
Vx5 xm5 0 0
Gx5_1 x5 0 u1 0 -0.0221441550850671
Rx6 x6 0 1
Fxc6_5 x6 0 Vx5 -8.7781784175362
Cx6 x6 xm6 1.3632937533957e-12
Vx6 xm6 0 0
Gx6_1 x6 0 u1 0 0.19438534424231
Rx7 x7 0 1
Fxc7_8 x7 0 Vx8 20.592055137168
Cx7 x7 xm7 6.0145717888717e-14
Vx7 xm7 0 0
Gx7_1 x7 0 u1 0 -0.000366486726882118
Rx8 x8 0 1
Fxc8_7 x8 0 Vx7 -4.17507177532355
Cx8 x8 xm8 6.0145717888717e-14
Vx8 xm8 0 0
Gx8_1 x8 0 u1 0 0.00153010838943624
Rx9 x9 0 1
Cx9 x9 0 7.61246317207855e-14
Gx9_1 x9 0 u1 0 -0.832460460165815
Rx10 x10 0 1
Cx10 x10 0 4.0771531282402e-13
Gx10_1 x10 0 u1 0 -1.77339574984073
Rx11 x11 0 1
Cx11 x11 0 3.62055457627861e-12
Gx11_1 x11 0 u1 0 -7.29153292860396
Rx12 x12 0 1
Fxc12_13 x12 0 Vx13 5.16250559123705
Cx12 x12 xm12 1.22121348511033e-13
Vx12 xm12 0 0
Gx12_2 x12 0 u2 0 -0.671027728999345
Rx13 x13 0 1
Fxc13_12 x13 0 Vx12 -0.632577257903099
Cx13 x13 xm13 1.22121348511033e-13
Vx13 xm13 0 0
Gx13_2 x13 0 u2 0 0.424476880787349
Rx14 x14 0 1
Fxc14_15 x14 0 Vx15 0.363608425840191
Cx14 x14 xm14 2.69558380066553e-12
Vx14 xm14 0 0
Gx14_2 x14 0 u2 0 -4.03228457762783
Rx15 x15 0 1
Fxc15_14 x15 0 Vx14 -0.372968257471828
Cx15 x15 xm15 2.69558380066553e-12
Vx15 xm15 0 0
Gx15_2 x15 0 u2 0 1.50391415254838
Rx16 x16 0 1
Fxc16_17 x16 0 Vx17 0.2825022999423
Cx16 x16 xm16 1.3632937533957e-12
Vx16 xm16 0 0
Gx16_2 x16 0 u2 0 -0.0205848577127193
Rx17 x17 0 1
Fxc17_16 x17 0 Vx16 -8.47001169799015
Cx17 x17 xm17 1.3632937533957e-12
Vx17 xm17 0 0
Gx17_2 x17 0 u2 0 0.174353985628195
Rx18 x18 0 1
Fxc18_19 x18 0 Vx19 13.9643157692737
Cx18 x18 xm18 6.0145717888717e-14
Vx18 xm18 0 0
Gx18_2 x18 0 u2 0 -0.000323685553711284
Rx19 x19 0 1
Fxc19_18 x19 0 Vx18 -6.15664309083206
Cx19 x19 xm19 6.0145717888717e-14
Vx19 xm19 0 0
Gx19_2 x19 0 u2 0 0.00199281642785873
Rx20 x20 0 1
Cx20 x20 0 7.61246317207855e-14
Gx20_2 x20 0 u2 0 -1.51377152400119
Rx21 x21 0 1
Cx21 x21 0 4.0771531282402e-13
Gx21_2 x21 0 u2 0 -1.77924060858146
Rx22 x22 0 1
Cx22 x22 0 3.62055457627861e-12
Gx22_2 x22 0 u2 0 -6.56797714514275
Gyc1_1 y1 0 x1 0 -0.435440967943983
Gyc1_2 y1 0 x2 0 1
Gyc1_3 y1 0 x3 0 1
Gyc1_4 y1 0 x4 0 -1
Gyc1_5 y1 0 x5 0 -1
Gyc1_6 y1 0 x6 0 1
Gyc1_7 y1 0 x7 0 1
Gyc1_8 y1 0 x8 0 -1
Gyc1_9 y1 0 x9 0 1
Gyc1_10 y1 0 x10 0 0.0922017921938196
Gyc1_11 y1 0 x11 0 -1
Gyc1_12 y1 0 x12 0 1
Gyc1_13 y1 0 x13 0 -0.156273052732549
Gyc1_14 y1 0 x14 0 -1
Gyc1_15 y1 0 x15 0 1
Gyc1_16 y1 0 x16 0 1
Gyc1_17 y1 0 x17 0 -1
Gyc1_18 y1 0 x18 0 -1
Gyc1_19 y1 0 x19 0 0.569209646365969
Gyc1_20 y1 0 x20 0 -0.137185636281771
Gyc1_21 y1 0 x21 0 -1
Gyc1_22 y1 0 x22 0 1
Gyc2_1 y2 0 x1 0 1
Gyc2_2 y2 0 x2 0 -0.199448689368593
Gyc2_3 y2 0 x3 0 -0.904004438616635
Gyc2_4 y2 0 x4 0 0.910598018472576
Gyc2_5 y2 0 x5 0 0.882269284478755
Gyc2_6 y2 0 x6 0 -0.90559082706608
Gyc2_7 y2 0 x7 0 -0.876870030643549
Gyc2_8 y2 0 x8 0 0.823325687673188
Gyc2_9 y2 0 x9 0 -0.253619876117991
Gyc2_10 y2 0 x10 0 -1
Gyc2_11 y2 0 x11 0 0.905730938531337
Gyc2_12 y2 0 x12 0 -0.980101215346374
Gyc2_13 y2 0 x13 0 -1
Gyc2_14 y2 0 x14 0 0.907982567043884
Gyc2_15 y2 0 x15 0 -0.933198535127717
Gyc2_16 y2 0 x16 0 -0.681423051117621
Gyc2_17 y2 0 x17 0 0.920682403656225
Gyc2_18 y2 0 x18 0 0.843049469132052
Gyc2_19 y2 0 x19 0 -1
Gyc2_20 y2 0 x20 0 1
Gyc2_21 y2 0 x21 0 -0.646859024742995
Gyc2_22 y2 0 x22 0 -0.913554325990294
.ENDS
