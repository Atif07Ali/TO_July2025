* Equivalent circuit model for E:\touchstone_files\inpmatch.ckt
.SUBCKT inpmatch po1 po2
Vsp1 po1 p1 0
Vsr1 p1 pr1 0
Rp1 pr1 0 50
Ru1 u1 0 50
Fr1 u1 0 Vsr1 -1
Fu1 u1 0 Vsp1 -1
Ry1 y1 0 1
Gy1 p1 0 y1 0 -0.02
Vsp2 po2 p2 0
Vsr2 p2 pr2 0
Rp2 pr2 0 50
Ru2 u2 0 50
Fr2 u2 0 Vsr2 -1
Fu2 u2 0 Vsp2 -1
Ry2 y2 0 1
Gy2 p2 0 y2 0 -0.02
Rx1 x1 0 1
Fxc1_2 x1 0 Vx2 12.3992364475181
Cx1 x1 xm1 1.44204939117694e-13
Vx1 xm1 0 0
Gx1_1 x1 0 u1 0 -0.606973349947336
Rx2 x2 0 1
Fxc2_1 x2 0 Vx1 -0.59924754498371
Cx2 x2 xm2 1.44204939117694e-13
Vx2 xm2 0 0
Gx2_1 x2 0 u1 0 0.363727289826479
Rx3 x3 0 1
Fxc3_4 x3 0 Vx4 3.95452200397614
Cx3 x3 xm3 2.6007985752599e-13
Vx3 xm3 0 0
Gx3_1 x3 0 u1 0 -0.496699864008767
Rx4 x4 0 1
Fxc4_3 x4 0 Vx3 -1.33880242756136
Cx4 x4 xm4 2.6007985752599e-13
Vx4 xm4 0 0
Gx4_1 x4 0 u1 0 0.664982983704334
Rx5 x5 0 1
Cx5 x5 0 1.16216062696842e-13
Gx5_1 x5 0 u1 0 -0.985547652963769
Rx6 x6 0 1
Cx6 x6 0 5.48902124943905e-13
Gx6_1 x6 0 u1 0 -1.44535589072413
Rx7 x7 0 1
Cx7 x7 0 3.80363316195477e-12
Gx7_1 x7 0 u1 0 -2.40718109029296
Rx8 x8 0 1
Fxc8_9 x8 0 Vx9 1.35052552994234
Cx8 x8 xm8 1.44204939117694e-13
Vx8 xm8 0 0
Gx8_2 x8 0 u2 0 -0.103484659623964
Rx9 x9 0 1
Fxc9_8 x9 0 Vx8 -5.50171902427121
Cx9 x9 xm9 1.44204939117694e-13
Vx9 xm9 0 0
Gx9_2 x9 0 u2 0 0.569343520573396
Rx10 x10 0 1
Fxc10_11 x10 0 Vx11 1.6536631180738
Cx10 x10 xm10 2.6007985752599e-13
Vx10 xm10 0 0
Gx10_2 x10 0 u2 0 -0.492390814796138
Rx11 x11 0 1
Fxc11_10 x11 0 Vx10 -3.20157328352036
Cx11 x11 xm11 2.6007985752599e-13
Vx11 xm11 0 0
Gx11_2 x11 0 u2 0 1.57642527770214
Rx12 x12 0 1
Cx12 x12 0 1.16216062696842e-13
Gx12_2 x12 0 u2 0 -0.880521652183412
Rx13 x13 0 1
Cx13 x13 0 5.48902124943906e-13
Gx13_2 x13 0 u2 0 -3.08436112780869
Rx14 x14 0 1
Cx14 x14 0 3.80363316195477e-12
Gx14_2 x14 0 u2 0 -0.833793414463596
Gyc1_1 y1 0 x1 0 -1
Gyc1_2 y1 0 x2 0 -0.838709870271279
Gyc1_3 y1 0 x3 0 -0.0940843337881672
Gyc1_4 y1 0 x4 0 1
Gyc1_5 y1 0 x5 0 1
Gyc1_6 y1 0 x6 0 1
Gyc1_7 y1 0 x7 0 -1
Gyc1_8 y1 0 x8 0 -1
Gyc1_9 y1 0 x9 0 0.620901184481792
Gyc1_10 y1 0 x10 0 1
Gyc1_11 y1 0 x11 0 0.308128194893076
Gyc1_12 y1 0 x12 0 -0.195347795861803
Gyc1_13 y1 0 x13 0 -0.0694754704557381
Gyc1_14 y1 0 x14 0 1
Gyc2_1 y2 0 x1 0 -0.178227780847756
Gyc2_2 y2 0 x2 0 1
Gyc2_3 y2 0 x3 0 1
Gyc2_4 y2 0 x4 0 0.781644854220982
Gyc2_5 y2 0 x5 0 -0.20622374645822
Gyc2_6 y2 0 x6 0 -0.0890649335462923
Gyc2_7 y2 0 x7 0 0.341670750101347
Gyc2_8 y2 0 x8 0 0.297127873334246
Gyc2_9 y2 0 x9 0 1
Gyc2_10 y2 0 x10 0 0.855308814147789
Gyc2_11 y2 0 x11 0 -1
Gyc2_12 y2 0 x12 0 1
Gyc2_13 y2 0 x13 0 -1
Gyc2_14 y2 0 x14 0 -0.29907384351315
.ENDS
