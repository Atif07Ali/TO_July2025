* Equivalent circuit model for E:\touchstone_files\output.ckt
.SUBCKT output po1 po2
Vsp1 po1 p1 0
Vsr1 p1 pr1 0
Rp1 pr1 0 50
Ru1 u1 0 50
Fr1 u1 0 Vsr1 -1
Fu1 u1 0 Vsp1 -1
Ry1 y1 0 1
Gy1 p1 0 y1 0 -0.02
Vsp2 po2 p2 0
Vsr2 p2 pr2 0
Rp2 pr2 0 50
Ru2 u2 0 50
Fr2 u2 0 Vsr2 -1
Fu2 u2 0 Vsp2 -1
Ry2 y2 0 1
Gy2 p2 0 y2 0 -0.02
Rx1 x1 0 1
Fxc1_2 x1 0 Vx2 2.19349705962773
Cx1 x1 xm1 2.97931551178328e-13
Vx1 xm1 0 0
Gx1_1 x1 0 u1 0 -0.774318205517317
Rx2 x2 0 1
Fxc2_1 x2 0 Vx1 -1.02146904001476
Cx2 x2 xm2 2.97931551178328e-13
Vx2 xm2 0 0
Gx2_1 x2 0 u1 0 0.790942074055725
Rx3 x3 0 1
Fxc3_4 x3 0 Vx4 7.90093857225456
Cx3 x3 xm3 5.60686590678349e-14
Vx3 xm3 0 0
Gx3_1 x3 0 u1 0 -0.121622272957677
Rx4 x4 0 1
Fxc4_3 x4 0 Vx3 -2.42192779343919
Cx4 x4 xm4 5.60686590678349e-14
Vx4 xm4 0 0
Gx4_1 x4 0 u1 0 0.294560363177445
Rx5 x5 0 1
Fxc5_6 x5 0 Vx6 7.33289855459071
Cx5 x5 xm5 2.36280354632591e-13
Vx5 xm5 0 0
Gx5_1 x5 0 u1 0 -0.0860988980115719
Rx6 x6 0 1
Fxc6_5 x6 0 Vx5 -1.86754985295544
Cx6 x6 xm6 2.36280354632591e-13
Vx6 xm6 0 0
Gx6_1 x6 0 u1 0 0.160793984321136
Rx7 x7 0 1
Fxc7_8 x7 0 Vx8 2.18178177801987
Cx7 x7 xm7 1.67762013258659e-13
Vx7 xm7 0 0
Gx7_1 x7 0 u1 0 -0.0230318402256142
Rx8 x8 0 1
Fxc8_7 x8 0 Vx7 -11.8287673323134
Cx8 x8 xm8 1.67762013258659e-13
Vx8 xm8 0 0
Gx8_1 x8 0 u1 0 0.272438279263806
Rx9 x9 0 1
Cx9 x9 0 9.66185966821205e-13
Gx9_1 x9 0 u1 0 -0.794072433112263
Rx10 x10 0 1
Fxc10_11 x10 0 Vx11 7.81833947606229
Cx10 x10 xm10 2.97931551178328e-13
Vx10 xm10 0 0
Gx10_2 x10 0 u2 0 -0.811122638261086
Rx11 x11 0 1
Fxc11_10 x11 0 Vx10 -0.286581228997952
Cx11 x11 xm11 2.97931551178328e-13
Vx11 xm11 0 0
Gx11_2 x11 0 u2 0 0.232452522540924
Rx12 x12 0 1
Fxc12_13 x12 0 Vx13 10.0036777508964
Cx12 x12 xm12 5.60686590678349e-14
Vx12 xm12 0 0
Gx12_2 x12 0 u2 0 -0.105674375595966
Rx13 x13 0 1
Fxc13_12 x13 0 Vx12 -1.91284677484583
Cx13 x13 xm13 5.6068659067835e-14
Vx13 xm13 0 0
Gx13_2 x13 0 u2 0 0.20213888854259
Rx14 x14 0 1
Fxc14_15 x14 0 Vx15 3.87902477535527
Cx14 x14 xm14 2.36280354632591e-13
Vx14 xm14 0 0
Gx14_2 x14 0 u2 0 -0.088307958249286
Rx15 x15 0 1
Fxc15_14 x15 0 Vx14 -3.53041148496113
Cx15 x15 xm15 2.36280354632591e-13
Vx15 xm15 0 0
Gx15_2 x15 0 u2 0 0.311763430016747
Rx16 x16 0 1
Fxc16_17 x16 0 Vx17 2.89649385601378
Cx16 x16 xm16 1.67762013258659e-13
Vx16 xm16 0 0
Gx16_2 x16 0 u2 0 -0.0331464746753219
Rx17 x17 0 1
Fxc17_16 x17 0 Vx16 -8.91000993097056
Cx17 x17 xm17 1.67762013258659e-13
Vx17 xm17 0 0
Gx17_2 x17 0 u2 0 0.295335418533782
Rx18 x18 0 1
Cx18 x18 0 9.66185966821205e-13
Gx18_2 x18 0 u2 0 -0.662072500089397
Gyc1_1 y1 0 x1 0 -0.262467472419468
Gyc1_2 y1 0 x2 0 -1
Gyc1_3 y1 0 x3 0 1
Gyc1_4 y1 0 x4 0 1
Gyc1_5 y1 0 x5 0 -1
Gyc1_6 y1 0 x6 0 0.909782426337428
Gyc1_7 y1 0 x7 0 -1
Gyc1_8 y1 0 x8 0 -0.075359970928032
Gyc1_9 y1 0 x9 0 1
Gyc1_10 y1 0 x10 0 -1
Gyc1_11 y1 0 x11 0 -0.330303290153262
Gyc1_12 y1 0 x12 0 1
Gyc1_13 y1 0 x13 0 -1
Gyc1_14 y1 0 x14 0 0.909649722032627
Gyc1_15 y1 0 x15 0 -0.659100474592723
Gyc1_16 y1 0 x16 0 1
Gyc1_17 y1 0 x17 0 -0.0273628799812312
Gyc1_18 y1 0 x18 0 0.147734907477295
Gyc2_1 y2 0 x1 0 -1
Gyc2_2 y2 0 x2 0 -0.360881176962411
Gyc2_3 y2 0 x3 0 0.871522390395498
Gyc2_4 y2 0 x4 0 -0.834509222992915
Gyc2_5 y2 0 x5 0 0.805215048233075
Gyc2_6 y2 0 x6 0 1
Gyc2_7 y2 0 x7 0 0.672947869535906
Gyc2_8 y2 0 x8 0 -1
Gyc2_9 y2 0 x9 0 -0.0768031605881768
Gyc2_10 y2 0 x10 0 0.189243483411446
Gyc2_11 y2 0 x11 0 -1
Gyc2_12 y2 0 x12 0 -0.213121763929887
Gyc2_13 y2 0 x13 0 -0.221368554324943
Gyc2_14 y2 0 x14 0 -1
Gyc2_15 y2 0 x15 0 -1
Gyc2_16 y2 0 x16 0 -0.703635239670564
Gyc2_17 y2 0 x17 0 1
Gyc2_18 y2 0 x18 0 1
.ENDS
