* Equivalent circuit model for E:\touchstone_files\interstage.ckt
.SUBCKT interstage po1 po2
Vsp1 po1 p1 0
Vsr1 p1 pr1 0
Rp1 pr1 0 50
Ru1 u1 0 50
Fr1 u1 0 Vsr1 -1
Fu1 u1 0 Vsp1 -1
Ry1 y1 0 1
Gy1 p1 0 y1 0 -0.02
Vsp2 po2 p2 0
Vsr2 p2 pr2 0
Rp2 pr2 0 50
Ru2 u2 0 50
Fr2 u2 0 Vsr2 -1
Fu2 u2 0 Vsp2 -1
Ry2 y2 0 1
Gy2 p2 0 y2 0 -0.02
Rx1 x1 0 1
Fxc1_2 x1 0 Vx2 0.786096295925692
Cx1 x1 xm1 2.20899391438717e-13
Vx1 xm1 0 0
Gx1_1 x1 0 u1 0 -0.540016668794603
Rx2 x2 0 1
Fxc2_1 x2 0 Vx1 -1.29688331062919
Cx2 x2 xm2 2.20899391438717e-13
Vx2 xm2 0 0
Gx2_1 x2 0 u1 0 0.700338605221292
Rx3 x3 0 1
Fxc3_4 x3 0 Vx4 19.6652440533082
Cx3 x3 xm3 9.54517955246503e-14
Vx3 xm3 0 0
Gx3_1 x3 0 u1 0 -0.0304277522431672
Rx4 x4 0 1
Fxc4_3 x4 0 Vx3 -2.50660661553957
Cx4 x4 xm4 9.54517955246503e-14
Vx4 xm4 0 0
Gx4_1 x4 0 u1 0 0.0762704050687221
Rx5 x5 0 1
Fxc5_6 x5 0 Vx6 26.2730628071917
Cx5 x5 xm5 7.14442889510699e-15
Vx5 xm5 0 0
Gx5_1 x5 0 u1 0 -4.26524034141191e-06
Rx6 x6 0 1
Fxc6_5 x6 0 Vx5 -458.728528471076
Cx6 x6 xm6 7.14442889510699e-15
Vx6 xm6 0 0
Gx6_1 x6 0 u1 0 0.00195658742539135
Rx7 x7 0 1
Fxc7_8 x7 0 Vx8 168.625431546935
Cx7 x7 xm7 2.94627305883564e-15
Vx7 xm7 0 0
Gx7_1 x7 0 u1 0 -1.19906563126763e-06
Rx8 x8 0 1
Fxc8_7 x8 0 Vx7 -208.739129538496
Cx8 x8 xm8 2.94627305883564e-15
Vx8 xm8 0 0
Gx8_1 x8 0 u1 0 0.000250291916130332
Rx9 x9 0 1
Cx9 x9 0 1.43904634962726e-12
Gx9_1 x9 0 u1 0 -1.2313168371131
Rx10 x10 0 1
Fxc10_11 x10 0 Vx11 1.00487572020899
Cx10 x10 xm10 2.20899391438717e-13
Vx10 xm10 0 0
Gx10_2 x10 0 u2 0 -0.646424214255343
Rx11 x11 0 1
Fxc11_10 x11 0 Vx10 -1.01452860909151
Cx11 x11 xm11 2.20899391438717e-13
Vx11 xm11 0 0
Gx11_2 x11 0 u2 0 0.655815858971543
Rx12 x12 0 1
Fxc12_13 x12 0 Vx13 34.9463368168507
Cx12 x12 xm12 9.54517955246503e-14
Vx12 xm12 0 0
Gx12_2 x12 0 u2 0 -0.0461848843997096
Rx13 x13 0 1
Fxc13_12 x13 0 Vx12 -1.41053498964888
Cx13 x13 xm13 9.54517955246503e-14
Vx13 xm13 0 0
Gx13_2 x13 0 u2 0 0.065145395438679
Rx14 x14 0 1
Fxc14_15 x14 0 Vx15 18.527826798324
Cx14 x14 xm14 7.14442889510699e-15
Vx14 xm14 0 0
Gx14_2 x14 0 u2 0 -4.18842128493827e-06
Rx15 x15 0 1
Fxc15_14 x15 0 Vx14 -650.492017825934
Cx15 x15 xm15 7.14442889510699e-15
Vx15 xm15 0 0
Gx15_2 x15 0 u2 0 0.00272453461314459
Rx16 x16 0 1
Fxc16_17 x16 0 Vx17 231.445889989574
Cx16 x16 xm16 2.94627305883564e-15
Vx16 xm16 0 0
Gx16_2 x16 0 u2 0 -2.74985141900546e-06
Rx17 x17 0 1
Fxc17_16 x17 0 Vx16 -152.08187883892
Cx17 x17 xm17 2.94627305883564e-15
Vx17 xm17 0 0
Gx17_2 x17 0 u2 0 0.000418202570330222
Rx18 x18 0 1
Cx18 x18 0 1.43904634962726e-12
Gx18_2 x18 0 u2 0 -1.22965625490186
Gyc1_1 y1 0 x1 0 1
Gyc1_2 y1 0 x2 0 -1
Gyc1_3 y1 0 x3 0 -0.653899698870499
Gyc1_4 y1 0 x4 0 1
Gyc1_5 y1 0 x5 0 0.979760723886354
Gyc1_6 y1 0 x6 0 0.77014328478896
Gyc1_7 y1 0 x7 0 -0.42232564894475
Gyc1_8 y1 0 x8 0 -0.0915503667380538
Gyc1_9 y1 0 x9 0 -0.931207271984113
Gyc1_10 y1 0 x10 0 0.0971351341549999
Gyc1_11 y1 0 x11 0 -0.111741261818517
Gyc1_12 y1 0 x12 0 0.659409096047566
Gyc1_13 y1 0 x13 0 -1
Gyc1_14 y1 0 x14 0 -1
Gyc1_15 y1 0 x15 0 -0.708237926203864
Gyc1_16 y1 0 x16 0 0.488004660046459
Gyc1_17 y1 0 x17 0 0.579286681215465
Gyc1_18 y1 0 x18 0 -1
Gyc2_1 y2 0 x1 0 0.110746723499143
Gyc2_2 y2 0 x2 0 -0.113857846865218
Gyc2_3 y2 0 x3 0 1
Gyc2_4 y2 0 x4 0 -0.82774151759558
Gyc2_5 y2 0 x5 0 -1
Gyc2_6 y2 0 x6 0 -1
Gyc2_7 y2 0 x7 0 1
Gyc2_8 y2 0 x8 0 1
Gyc2_9 y2 0 x9 0 -1
Gyc2_10 y2 0 x10 0 1
Gyc2_11 y2 0 x11 0 -1
Gyc2_12 y2 0 x12 0 -1
Gyc2_13 y2 0 x13 0 0.559911956021983
Gyc2_14 y2 0 x14 0 0.847318039595005
Gyc2_15 y2 0 x15 0 1
Gyc2_16 y2 0 x16 0 -1
Gyc2_17 y2 0 x17 0 -1
Gyc2_18 y2 0 x18 0 -0.992739409346559
.ENDS
