* Equivalent circuit model for E:\touchstone_files\choke_last5.s3p.ckt
.SUBCKT choke_last5.s3p po1 po2 po3
Vsp1 po1 p1 0
Vsr1 p1 pr1 0
Rp1 pr1 0 50
Ru1 u1 0 50
Fr1 u1 0 Vsr1 -1
Fu1 u1 0 Vsp1 -1
Ry1 y1 0 1
Gy1 p1 0 y1 0 -0.02
Vsp2 po2 p2 0
Vsr2 p2 pr2 0
Rp2 pr2 0 50
Ru2 u2 0 50
Fr2 u2 0 Vsr2 -1
Fu2 u2 0 Vsp2 -1
Ry2 y2 0 1
Gy2 p2 0 y2 0 -0.02
Vsp3 po3 p3 0
Vsr3 p3 pr3 0
Rp3 pr3 0 50
Ru3 u3 0 50
Fr3 u3 0 Vsr3 -1
Fu3 u3 0 Vsp3 -1
Ry3 y3 0 1
Gy3 p3 0 y3 0 -0.02
Rx1 x1 0 1
Fxc1_2 x1 0 Vx2 1.77205808235061
Cx1 x1 xm1 1.43937031105238e-13
Vx1 xm1 0 0
Gx1_1 x1 0 u1 0 -0.109979031423695
Rx2 x2 0 1
Fxc2_1 x2 0 Vx1 -4.80049636089305
Cx2 x2 xm2 1.43937031105238e-13
Vx2 xm2 0 0
Gx2_1 x2 0 u1 0 0.527953940123991
Rx3 x3 0 1
Fxc3_4 x3 0 Vx4 0.385547237492729
Cx3 x3 xm3 5.71274901965996e-13
Vx3 xm3 0 0
Gx3_1 x3 0 u1 0 -0.163082001364491
Rx4 x4 0 1
Fxc4_3 x4 0 Vx3 -3.91600491344283
Cx4 x4 xm4 5.71274901965996e-13
Vx4 xm4 0 0
Gx4_1 x4 0 u1 0 0.638629918637435
Rx5 x5 0 1
Fxc5_6 x5 0 Vx6 6.60657201620162
Cx5 x5 xm5 2.40075948885019e-13
Vx5 xm5 0 0
Gx5_1 x5 0 u1 0 -0.0255787526861871
Rx6 x6 0 1
Fxc6_5 x6 0 Vx5 -2.55607599735171
Cx6 x6 xm6 2.40075948885019e-13
Vx6 xm6 0 0
Gx6_1 x6 0 u1 0 0.0653812357833583
Rx7 x7 0 1
Fxc7_8 x7 0 Vx8 1.67988510588745
Cx7 x7 xm7 6.05230657216695e-14
Vx7 xm7 0 0
Gx7_1 x7 0 u1 0 -0.00219539790391067
Rx8 x8 0 1
Fxc8_7 x8 0 Vx7 -52.7646908890623
Cx8 x8 xm8 6.05230657216695e-14
Vx8 xm8 0 0
Gx8_1 x8 0 u1 0 0.115839491778342
Rx9 x9 0 1
Fxc9_10 x9 0 Vx10 0.763692255550998
Cx9 x9 xm9 4.41970619749814e-12
Vx9 xm9 0 0
Gx9_1 x9 0 u1 0 -2.57870099673024
Rx10 x10 0 1
Fxc10_9 x10 0 Vx9 -0.615819680772403
Cx10 x10 xm10 4.41970619749814e-12
Vx10 xm10 0 0
Gx10_1 x10 0 u1 0 1.58801482461389
Rx11 x11 0 1
Fxc11_12 x11 0 Vx12 5.9074668073064
Cx11 x11 xm11 2.20312369841031e-12
Vx11 xm11 0 0
Gx11_1 x11 0 u1 0 -1.49895091570117
Rx12 x12 0 1
Fxc12_11 x12 0 Vx11 -0.41402306443572
Cx12 x12 xm12 2.20312369841031e-12
Vx12 xm12 0 0
Gx12_1 x12 0 u1 0 0.620600251557327
Rx13 x13 0 1
Fxc13_14 x13 0 Vx14 3.175223871049
Cx13 x13 xm13 4.22338545561999e-14
Vx13 xm13 0 0
Gx13_1 x13 0 u1 0 -0.000782184042617225
Rx14 x14 0 1
Fxc14_13 x14 0 Vx13 -59.9039123466464
Cx14 x14 xm14 4.22338545561999e-14
Vx14 xm14 0 0
Gx14_1 x14 0 u1 0 0.0468558843278878
Rx15 x15 0 1
Fxc15_16 x15 0 Vx16 0.200069031213313
Cx15 x15 xm15 8.2912818041689e-13
Vx15 xm15 0 0
Gx15_1 x15 0 u1 0 -0.00511150073777445
Rx16 x16 0 1
Fxc16_15 x16 0 Vx15 -55.0120979235847
Cx16 x16 xm16 8.2912818041689e-13
Vx16 xm16 0 0
Gx16_1 x16 0 u1 0 0.281194379122923
Rx17 x17 0 1
Fxc17_18 x17 0 Vx18 15.6957310166792
Cx17 x17 xm17 3.97491807667442e-14
Vx17 xm17 0 0
Gx17_1 x17 0 u1 0 -0.000281806144110906
Rx18 x18 0 1
Fxc18_17 x18 0 Vx17 -16.6821734613482
Cx18 x18 xm18 3.97491807667442e-14
Vx18 xm18 0 0
Gx18_1 x18 0 u1 0 0.00470113897853184
Rx19 x19 0 1
Fxc19_20 x19 0 Vx20 26.5067987561139
Cx19 x19 xm19 2.48712484007818e-14
Vx19 xm19 0 0
Gx19_1 x19 0 u1 0 -0.000404733917101592
Rx20 x20 0 1
Fxc20_19 x20 0 Vx19 -17.4975920781252
Cx20 x20 xm20 2.48712484007818e-14
Vx20 xm20 0 0
Gx20_1 x20 0 u1 0 0.00708186898162538
Rx21 x21 0 1
Fxc21_22 x21 0 Vx22 2.71365477347699
Cx21 x21 xm21 2.87619707206074e-13
Vx21 xm21 0 0
Gx21_1 x21 0 u1 0 -0.00120530358282358
Rx22 x22 0 1
Fxc22_21 x22 0 Vx21 -17.4614505440889
Cx22 x22 xm22 2.87619707206074e-13
Vx22 xm22 0 0
Gx22_1 x22 0 u1 0 0.0210463489020871
Rx23 x23 0 1
Fxc23_24 x23 0 Vx24 10.119964335474
Cx23 x23 xm23 3.56268627400195e-14
Vx23 xm23 0 0
Gx23_1 x23 0 u1 0 -2.74077954554101e-05
Rx24 x24 0 1
Fxc24_23 x24 0 Vx23 -45.1574490319763
Cx24 x24 xm24 3.56268627400195e-14
Vx24 xm24 0 0
Gx24_1 x24 0 u1 0 0.00123766612635651
Rx25 x25 0 1
Fxc25_26 x25 0 Vx26 42.6011900965731
Cx25 x25 xm25 1.2637138685889e-13
Vx25 xm25 0 0
Gx25_1 x25 0 u1 0 -0.000362421654159091
Rx26 x26 0 1
Fxc26_25 x26 0 Vx25 -3.13721196943335
Cx26 x26 xm26 1.2637138685889e-13
Vx26 xm26 0 0
Gx26_1 x26 0 u1 0 0.00113699355140973
Rx27 x27 0 1
Cx27 x27 0 7.65184566999521e-12
Gx27_1 x27 0 u1 0 -1.30069142311978
Rx28 x28 0 1
Fxc28_29 x28 0 Vx29 1.40263720560015
Cx28 x28 xm28 1.43937031105238e-13
Vx28 xm28 0 0
Gx28_2 x28 0 u2 0 -0.0980870979251834
Rx29 x29 0 1
Fxc29_28 x29 0 Vx28 -6.06483154849396
Cx29 x29 xm29 1.43937031105238e-13
Vx29 xm29 0 0
Gx29_2 x29 0 u2 0 0.594881725996869
Rx30 x30 0 1
Fxc30_31 x30 0 Vx31 0.606513445551286
Cx30 x30 xm30 5.71274901965996e-13
Vx30 xm30 0 0
Gx30_2 x30 0 u2 0 -0.232297858324788
Rx31 x31 0 1
Fxc31_30 x31 0 Vx30 -2.48931806452124
Cx31 x31 xm31 5.71274901965996e-13
Vx31 xm31 0 0
Gx31_2 x31 0 u2 0 0.578263255077491
Rx32 x32 0 1
Fxc32_33 x32 0 Vx33 2.68120549956711
Cx32 x32 xm32 2.40075948885019e-13
Vx32 xm32 0 0
Gx32_2 x32 0 u2 0 -0.0168679139035021
Rx33 x33 0 1
Fxc33_32 x33 0 Vx32 -6.29824911149665
Cx33 x33 xm33 2.40075948885019e-13
Vx33 xm33 0 0
Gx33_2 x33 0 u2 0 0.106238323755534
Rx34 x34 0 1
Fxc34_35 x34 0 Vx35 8.1458023300897
Cx34 x34 xm34 6.05230657216695e-14
Vx34 xm34 0 0
Gx34_2 x34 0 u2 0 -0.00993474379877102
Rx35 x35 0 1
Fxc35_34 x35 0 Vx34 -10.8815086285448
Cx35 x35 xm35 6.05230657216695e-14
Vx35 xm35 0 0
Gx35_2 x35 0 u2 0 0.108105000368709
Rx36 x36 0 1
Fxc36_37 x36 0 Vx37 0.911839983568162
Cx36 x36 xm36 4.41970619749814e-12
Vx36 xm36 0 0
Gx36_2 x36 0 u2 0 -2.8639587646356
Rx37 x37 0 1
Fxc37_36 x37 0 Vx36 -0.515766723873451
Cx37 x37 xm37 4.41970619749814e-12
Vx37 xm37 0 0
Gx37_2 x37 0 u2 0 1.47713462934476
Rx38 x38 0 1
Fxc38_39 x38 0 Vx39 3.32650853258027
Cx38 x38 xm38 2.20312369841031e-12
Vx38 xm38 0 0
Gx38_2 x38 0 u2 0 -1.49839134997013
Rx39 x39 0 1
Fxc39_38 x39 0 Vx38 -0.735253641064957
Cx39 x39 xm39 2.20312369841031e-12
Vx39 xm39 0 0
Gx39_2 x39 0 u2 0 1.10169769580578
Rx40 x40 0 1
Fxc40_41 x40 0 Vx41 8.15973187889306
Cx40 x40 xm40 4.22338545561999e-14
Vx40 xm40 0 0
Gx40_2 x40 0 u2 0 -0.0020641677267741
Rx41 x41 0 1
Fxc41_40 x41 0 Vx40 -23.3106106028207
Cx41 x41 xm41 4.22338545561999e-14
Vx41 xm41 0 0
Gx41_2 x41 0 u2 0 0.0481170100977406
Rx42 x42 0 1
Fxc42_43 x42 0 Vx43 0.739187322844793
Cx42 x42 xm42 8.2912818041689e-13
Vx42 xm42 0 0
Gx42_2 x42 0 u2 0 -0.0191731559373127
Rx43 x43 0 1
Fxc43_42 x43 0 Vx42 -14.8896183638886
Cx43 x43 xm43 8.2912818041689e-13
Vx43 xm43 0 0
Gx43_2 x43 0 u2 0 0.285480974737911
Rx44 x44 0 1
Fxc44_45 x44 0 Vx45 4.36026229800473
Cx44 x44 xm44 3.97491807667442e-14
Vx44 xm44 0 0
Gx44_2 x44 0 u2 0 -0.000107433314512435
Rx45 x45 0 1
Fxc45_44 x45 0 Vx44 -60.0511825957638
Cx45 x45 xm45 3.97491807667442e-14
Vx45 xm45 0 0
Gx45_2 x45 0 u2 0 0.00645149758665435
Rx46 x46 0 1
Fxc46_47 x46 0 Vx47 279.288761629974
Cx46 x46 xm46 2.48712484007818e-14
Vx46 xm46 0 0
Gx46_2 x46 0 u2 0 -0.000581160552840632
Rx47 x47 0 1
Fxc47_46 x47 0 Vx46 -1.66066528858733
Cx47 x47 xm47 2.48712484007818e-14
Vx47 xm47 0 0
Gx47_2 x47 0 u2 0 0.000965113157198657
Rx48 x48 0 1
Fxc48_49 x48 0 Vx49 3.98363562554835
Cx48 x48 xm48 2.87619707206074e-13
Vx48 xm48 0 0
Gx48_2 x48 0 u2 0 -0.00163464550223602
Rx49 x49 0 1
Fxc49_48 x49 0 Vx48 -11.8947496896825
Cx49 x49 xm49 2.87619707206074e-13
Vx49 xm49 0 0
Gx49_2 x49 0 u2 0 0.0194436990804628
Rx50 x50 0 1
Fxc50_51 x50 0 Vx51 8.71705145459893
Cx50 x50 xm50 3.56268627400195e-14
Vx50 xm50 0 0
Gx50_2 x50 0 u2 0 -1.94929483067017e-05
Rx51 x51 0 1
Fxc51_50 x51 0 Vx50 -52.425040286241
Cx51 x51 xm51 3.56268627400195e-14
Vx51 xm51 0 0
Gx51_2 x51 0 u2 0 0.00102191860027645
Rx52 x52 0 1
Fxc52_53 x52 0 Vx53 23.1337493790108
Cx52 x52 xm52 1.2637138685889e-13
Vx52 xm52 0 0
Gx52_2 x52 0 u2 0 -0.000323078412656316
Rx53 x53 0 1
Fxc53_52 x53 0 Vx52 -5.77722881377516
Cx53 x53 xm53 1.2637138685889e-13
Vx53 xm53 0 0
Gx53_2 x53 0 u2 0 0.00186649791470681
Rx54 x54 0 1
Cx54 x54 0 7.65184566999521e-12
Gx54_2 x54 0 u2 0 -1.65787522447043
Rx55 x55 0 1
Fxc55_56 x55 0 Vx56 77.8534997478518
Cx55 x55 xm55 1.43937031105238e-13
Vx55 xm55 0 0
Gx55_3 x55 0 u3 0 -0.662441964373491
Rx56 x56 0 1
Fxc56_55 x56 0 Vx55 -0.109266229561503
Cx56 x56 xm56 1.43937031105238e-13
Vx56 xm56 0 0
Gx56_3 x56 0 u3 0 0.0723825357504071
Rx57 x57 0 1
Fxc57_58 x57 0 Vx58 2.23171058279709
Cx57 x57 xm57 5.71274901965996e-13
Vx57 xm57 0 0
Gx57_3 x57 0 u3 0 -4.52124469300687
Rx58 x58 0 1
Fxc58_57 x58 0 Vx57 -0.676523599441618
Cx58 x58 xm58 5.71274901965996e-13
Vx58 xm58 0 0
Gx58_3 x58 0 u3 0 3.05872873366932
Rx59 x59 0 1
Fxc59_60 x59 0 Vx60 93.4449409487633
Cx59 x59 xm59 2.40075948885019e-13
Vx59 xm59 0 0
Gx59_3 x59 0 u3 0 -0.500337113727103
Rx60 x60 0 1
Fxc60_59 x60 0 Vx59 -0.180714974871114
Cx60 x60 xm60 2.40075948885019e-13
Vx60 xm60 0 0
Gx60_3 x60 0 u3 0 0.090418408934279
Rx61 x61 0 1
Fxc61_62 x61 0 Vx62 2.2772994665264
Cx61 x61 xm61 6.05230657216695e-14
Vx61 xm61 0 0
Gx61_3 x61 0 u3 0 -0.0145915097577578
Rx62 x62 0 1
Fxc62_61 x62 0 Vx61 -38.9226887566496
Cx62 x62 xm62 6.05230657216695e-14
Vx62 xm62 0 0
Gx62_3 x62 0 u3 0 0.567940792790823
Rx63 x63 0 1
Fxc63_64 x63 0 Vx64 0.678695999944544
Cx63 x63 xm63 4.41970619749814e-12
Vx63 xm63 0 0
Gx63_3 x63 0 u3 0 -2.06450091695134
Rx64 x64 0 1
Fxc64_63 x64 0 Vx63 -0.692941642591381
Cx64 x64 xm64 4.41970619749814e-12
Vx64 xm64 0 0
Gx64_3 x64 0 u3 0 1.43057865652368
Rx65 x65 0 1
Fxc65_66 x65 0 Vx66 2.25797191566121
Cx65 x65 xm65 2.20312369841031e-12
Vx65 xm65 0 0
Gx65_3 x65 0 u3 0 -0.700618752856902
Rx66 x66 0 1
Fxc66_65 x66 0 Vx65 -1.08319660384132
Cx66 x66 xm66 2.20312369841031e-12
Vx66 xm66 0 0
Gx66_3 x66 0 u3 0 0.758907853682135
Rx67 x67 0 1
Fxc67_68 x67 0 Vx68 18.4679823140632
Cx67 x67 xm67 4.22338545561999e-14
Vx67 xm67 0 0
Gx67_3 x67 0 u3 0 -0.00482038020061546
Rx68 x68 0 1
Fxc68_67 x68 0 Vx67 -10.2993564330769
Cx68 x68 xm68 4.22338545561998e-14
Vx68 xm68 0 0
Gx68_3 x68 0 u3 0 0.0496468138290856
Rx69 x69 0 1
Fxc69_70 x69 0 Vx70 5.94381439194125
Cx69 x69 xm69 8.2912818041689e-13
Vx69 xm69 0 0
Gx69_3 x69 0 u3 0 -0.0329355480014432
Rx70 x70 0 1
Fxc70_69 x70 0 Vx69 -1.85170942610623
Cx70 x70 xm70 8.2912818041689e-13
Vx70 xm70 0 0
Gx70_3 x70 0 u3 0 0.0609870646882466
Rx71 x71 0 1
Fxc71_72 x71 0 Vx72 129.471905479814
Cx71 x71 xm71 3.97491807667442e-14
Vx71 xm71 0 0
Gx71_3 x71 0 u3 0 -0.000934132271612798
Rx72 x72 0 1
Fxc72_71 x72 0 Vx71 -2.0223608083356
Cx72 x72 xm72 3.97491807667442e-14
Vx72 xm72 0 0
Gx72_3 x72 0 u3 0 0.00188915249591123
Rx73 x73 0 1
Fxc73_74 x73 0 Vx74 71.4001954230967
Cx73 x73 xm73 2.48712484007818e-14
Vx73 xm73 0 0
Gx73_3 x73 0 u3 0 -0.00029563792428037
Rx74 x74 0 1
Fxc74_73 x74 0 Vx73 -6.4958526959634
Cx74 x74 xm74 2.48712484007817e-14
Vx74 xm74 0 0
Gx74_3 x74 0 u3 0 0.00192042040746566
Rx75 x75 0 1
Fxc75_76 x75 0 Vx76 12.5648465121659
Cx75 x75 xm75 2.87619707206074e-13
Vx75 xm75 0 0
Gx75_3 x75 0 u3 0 -0.00122687327540189
Rx76 x76 0 1
Fxc76_75 x76 0 Vx75 -3.77118403913009
Cx76 x76 xm76 2.87619707206074e-13
Vx76 xm76 0 0
Gx76_3 x76 0 u3 0 0.00462676491423088
Rx77 x77 0 1
Fxc77_78 x77 0 Vx78 18.7097601595856
Cx77 x77 xm77 3.56268627400195e-14
Vx77 xm77 0 0
Gx77_3 x77 0 u3 0 -0.00011756152141632
Rx78 x78 0 1
Fxc78_77 x78 0 Vx77 -24.4253143699682
Cx78 x78 xm78 3.56268627400195e-14
Vx78 xm78 0 0
Gx78_3 x78 0 u3 0 0.00287147711840536
Rx79 x79 0 1
Fxc79_80 x79 0 Vx80 17.0697363591418
Cx79 x79 xm79 1.2637138685889e-13
Vx79 xm79 0 0
Gx79_3 x79 0 u3 0 -0.000144706394217082
Rx80 x80 0 1
Fxc80_79 x80 0 Vx79 -7.82958568727381
Cx80 x80 xm80 1.2637138685889e-13
Vx80 xm80 0 0
Gx80_3 x80 0 u3 0 0.00113299111301907
Rx81 x81 0 1
Cx81 x81 0 7.65184566999521e-12
Gx81_3 x81 0 u3 0 -2.35910769694722
Gyc1_1 y1 0 x1 0 -1
Gyc1_2 y1 0 x2 0 -1
Gyc1_3 y1 0 x3 0 0.203839141557435
Gyc1_4 y1 0 x4 0 -1
Gyc1_5 y1 0 x5 0 0.212149977103385
Gyc1_6 y1 0 x6 0 0.633843378159311
Gyc1_7 y1 0 x7 0 -1
Gyc1_8 y1 0 x8 0 -0.613728845299851
Gyc1_9 y1 0 x9 0 1
Gyc1_10 y1 0 x10 0 1
Gyc1_11 y1 0 x11 0 -1
Gyc1_12 y1 0 x12 0 0.885533835328313
Gyc1_13 y1 0 x13 0 -0.201437357973855
Gyc1_14 y1 0 x14 0 0.768409848201219
Gyc1_15 y1 0 x15 0 0.0629452490909661
Gyc1_16 y1 0 x16 0 -0.944534278392737
Gyc1_17 y1 0 x17 0 -0.78669079814722
Gyc1_18 y1 0 x18 0 1
Gyc1_19 y1 0 x19 0 0.549996341374664
Gyc1_20 y1 0 x20 0 1
Gyc1_21 y1 0 x21 0 -0.718554247020533
Gyc1_22 y1 0 x22 0 -0.959243997194098
Gyc1_23 y1 0 x23 0 0.0155509826328834
Gyc1_24 y1 0 x24 0 -1
Gyc1_25 y1 0 x25 0 -1
Gyc1_26 y1 0 x26 0 0.580503341865985
Gyc1_27 y1 0 x27 0 -0.0153977387617627
Gyc1_28 y1 0 x28 0 -0.512953194423879
Gyc1_29 y1 0 x29 0 0.0628197106145299
Gyc1_30 y1 0 x30 0 1
Gyc1_31 y1 0 x31 0 0.384443465745625
Gyc1_32 y1 0 x32 0 -0.381035709132174
Gyc1_33 y1 0 x33 0 -0.101125739794263
Gyc1_34 y1 0 x34 0 0.773104759911681
Gyc1_35 y1 0 x35 0 1
Gyc1_36 y1 0 x36 0 -0.773968267076957
Gyc1_37 y1 0 x37 0 -1
Gyc1_38 y1 0 x38 0 1
Gyc1_39 y1 0 x39 0 -0.628037874188683
Gyc1_40 y1 0 x40 0 -0.681963105850894
Gyc1_41 y1 0 x41 0 -1
Gyc1_42 y1 0 x42 0 0.591801771193975
Gyc1_43 y1 0 x43 0 1
Gyc1_44 y1 0 x44 0 1
Gyc1_45 y1 0 x45 0 -0.934649292141004
Gyc1_46 y1 0 x46 0 -1
Gyc1_47 y1 0 x47 0 1
Gyc1_48 y1 0 x48 0 1
Gyc1_49 y1 0 x49 0 1
Gyc1_50 y1 0 x50 0 0.721298725674352
Gyc1_51 y1 0 x51 0 0.929270107184347
Gyc1_52 y1 0 x52 0 1
Gyc1_53 y1 0 x53 0 -1
Gyc1_54 y1 0 x54 0 -1
Gyc1_55 y1 0 x55 0 -0.0417301419330315
Gyc1_56 y1 0 x56 0 -0.0239498126563669
Gyc1_57 y1 0 x57 0 0.032160235415803
Gyc1_58 y1 0 x58 0 0.0872445937942062
Gyc1_59 y1 0 x59 0 -0.0546072574008846
Gyc1_60 y1 0 x60 0 -1
Gyc1_61 y1 0 x61 0 -0.108908376302564
Gyc1_62 y1 0 x62 0 0.0723608705676596
Gyc1_63 y1 0 x63 0 1
Gyc1_64 y1 0 x64 0 0.853963280804006
Gyc1_65 y1 0 x65 0 -0.954977821009915
Gyc1_66 y1 0 x66 0 0.995069370846795
Gyc1_67 y1 0 x67 0 0.0808136288042712
Gyc1_68 y1 0 x68 0 -0.263516160347489
Gyc1_69 y1 0 x69 0 -0.813198071595963
Gyc1_70 y1 0 x70 0 -0.866282997260543
Gyc1_71 y1 0 x71 0 0.193488735789555
Gyc1_72 y1 0 x72 0 -0.514146022555978
Gyc1_73 y1 0 x73 0 -0.428040729744565
Gyc1_74 y1 0 x74 0 -0.2261853293714
Gyc1_75 y1 0 x75 0 -0.697503489687245
Gyc1_76 y1 0 x76 0 0.6328360512145
Gyc1_77 y1 0 x77 0 0.0829238674504882
Gyc1_78 y1 0 x78 0 0.158305795298448
Gyc1_79 y1 0 x79 0 0.457555141700982
Gyc1_80 y1 0 x80 0 0.560513607129299
Gyc1_81 y1 0 x81 0 0.00958620036356174
Gyc2_1 y2 0 x1 0 -0.327792642991468
Gyc2_2 y2 0 x2 0 -0.0365945474106578
Gyc2_3 y2 0 x3 0 1
Gyc2_4 y2 0 x4 0 0.411589821142152
Gyc2_5 y2 0 x5 0 -0.192610490353332
Gyc2_6 y2 0 x6 0 -0.270261566592714
Gyc2_7 y2 0 x7 0 -0.0518401785495051
Gyc2_8 y2 0 x8 0 1
Gyc2_9 y2 0 x9 0 -0.777564305386856
Gyc2_10 y2 0 x10 0 -0.71094011042537
Gyc2_11 y2 0 x11 0 0.933339290074078
Gyc2_12 y2 0 x12 0 -1
Gyc2_13 y2 0 x13 0 1
Gyc2_14 y2 0 x14 0 -1
Gyc2_15 y2 0 x15 0 0.700070261033951
Gyc2_16 y2 0 x16 0 1
Gyc2_17 y2 0 x17 0 1
Gyc2_18 y2 0 x18 0 -0.896414537811581
Gyc2_19 y2 0 x19 0 -1
Gyc2_20 y2 0 x20 0 -0.932055584476272
Gyc2_21 y2 0 x21 0 1
Gyc2_22 y2 0 x22 0 1
Gyc2_23 y2 0 x23 0 -0.247561313615287
Gyc2_24 y2 0 x24 0 0.8360379689621
Gyc2_25 y2 0 x25 0 0.989313295789868
Gyc2_26 y2 0 x26 0 -1
Gyc2_27 y2 0 x27 0 -1
Gyc2_28 y2 0 x28 0 -1
Gyc2_29 y2 0 x29 0 -1
Gyc2_30 y2 0 x30 0 -0.136701603627477
Gyc2_31 y2 0 x31 0 -1
Gyc2_32 y2 0 x32 0 0.31326107186107
Gyc2_33 y2 0 x33 0 0.294158767613144
Gyc2_34 y2 0 x34 0 -1
Gyc2_35 y2 0 x35 0 -0.513407195759489
Gyc2_36 y2 0 x36 0 1
Gyc2_37 y2 0 x37 0 0.695990582752553
Gyc2_38 y2 0 x38 0 -0.920167170720914
Gyc2_39 y2 0 x39 0 1
Gyc2_40 y2 0 x40 0 1
Gyc2_41 y2 0 x41 0 0.718001787486554
Gyc2_42 y2 0 x42 0 -1
Gyc2_43 y2 0 x43 0 -0.904814247463402
Gyc2_44 y2 0 x44 0 -0.253706250212905
Gyc2_45 y2 0 x45 0 1
Gyc2_46 y2 0 x46 0 0.615351651468943
Gyc2_47 y2 0 x47 0 -0.540962676315279
Gyc2_48 y2 0 x48 0 -0.93053255686352
Gyc2_49 y2 0 x49 0 -0.902186906579574
Gyc2_50 y2 0 x50 0 -1
Gyc2_51 y2 0 x51 0 -1
Gyc2_52 y2 0 x52 0 -0.991322318920966
Gyc2_53 y2 0 x53 0 0.828936290595289
Gyc2_54 y2 0 x54 0 -0.223494342321579
Gyc2_55 y2 0 x55 0 0.0516243139048618
Gyc2_56 y2 0 x56 0 0.184340089189232
Gyc2_57 y2 0 x57 0 0.00579588735582951
Gyc2_58 y2 0 x58 0 -0.111042047790681
Gyc2_59 y2 0 x59 0 -0.0296224922305034
Gyc2_60 y2 0 x60 0 -0.844022815342035
Gyc2_61 y2 0 x61 0 0.209901768540489
Gyc2_62 y2 0 x62 0 -0.0982392171106038
Gyc2_63 y2 0 x63 0 -0.797804308001655
Gyc2_64 y2 0 x64 0 -1
Gyc2_65 y2 0 x65 0 1
Gyc2_66 y2 0 x66 0 -1
Gyc2_67 y2 0 x67 0 -0.18419063456975
Gyc2_68 y2 0 x68 0 0.283830335675255
Gyc2_69 y2 0 x69 0 1
Gyc2_70 y2 0 x70 0 1
Gyc2_71 y2 0 x71 0 -0.196870786594296
Gyc2_72 y2 0 x72 0 0.168121850202167
Gyc2_73 y2 0 x73 0 0.459694579026774
Gyc2_74 y2 0 x74 0 1
Gyc2_75 y2 0 x75 0 1
Gyc2_76 y2 0 x76 0 -1
Gyc2_77 y2 0 x77 0 0.16972702074558
Gyc2_78 y2 0 x78 0 -0.200672217220817
Gyc2_79 y2 0 x79 0 -1
Gyc2_80 y2 0 x80 0 -1
Gyc2_81 y2 0 x81 0 -1
Gyc3_1 y3 0 x1 0 0.0768182204483113
Gyc3_2 y3 0 x2 0 -0.000669197600108597
Gyc3_3 y3 0 x3 0 0.494349856480557
Gyc3_4 y3 0 x4 0 -0.121436726891915
Gyc3_5 y3 0 x5 0 -1
Gyc3_6 y3 0 x6 0 -1
Gyc3_7 y3 0 x7 0 -0.570160867535789
Gyc3_8 y3 0 x8 0 -0.214810827156227
Gyc3_9 y3 0 x9 0 0.450008577977847
Gyc3_10 y3 0 x10 0 0.133320099016962
Gyc3_11 y3 0 x11 0 -0.283418456453302
Gyc3_12 y3 0 x12 0 0.662636652333409
Gyc3_13 y3 0 x13 0 -0.311783848314679
Gyc3_14 y3 0 x14 0 0.221212502657933
Gyc3_15 y3 0 x15 0 -1
Gyc3_16 y3 0 x16 0 -0.26802616178998
Gyc3_17 y3 0 x17 0 -0.143745397086877
Gyc3_18 y3 0 x18 0 0.0759293707485176
Gyc3_19 y3 0 x19 0 0.192680897466469
Gyc3_20 y3 0 x20 0 0.2027179721114
Gyc3_21 y3 0 x21 0 -0.235302408210299
Gyc3_22 y3 0 x22 0 -0.261614704266111
Gyc3_23 y3 0 x23 0 1
Gyc3_24 y3 0 x24 0 -0.278857416644056
Gyc3_25 y3 0 x25 0 -0.3225868303356
Gyc3_26 y3 0 x26 0 0.0293780559531698
Gyc3_27 y3 0 x27 0 -0.821501605888946
Gyc3_28 y3 0 x28 0 -0.146180802210975
Gyc3_29 y3 0 x29 0 0.0258625412226248
Gyc3_30 y3 0 x30 0 0.489824504478502
Gyc3_31 y3 0 x31 0 0.169553664895352
Gyc3_32 y3 0 x32 0 -1
Gyc3_33 y3 0 x33 0 -1
Gyc3_34 y3 0 x34 0 0.422689399999568
Gyc3_35 y3 0 x35 0 0.297395427720841
Gyc3_36 y3 0 x36 0 -0.178589680146573
Gyc3_37 y3 0 x37 0 -0.14309748579302
Gyc3_38 y3 0 x38 0 0.273723533954663
Gyc3_39 y3 0 x39 0 -0.291367868461571
Gyc3_40 y3 0 x40 0 -0.26336084760432
Gyc3_41 y3 0 x41 0 -0.383316117511786
Gyc3_42 y3 0 x42 0 0.357762872972679
Gyc3_43 y3 0 x43 0 0.329898007484434
Gyc3_44 y3 0 x44 0 0.467134282132148
Gyc3_45 y3 0 x45 0 -0.306214024806134
Gyc3_46 y3 0 x46 0 -0.34374591936894
Gyc3_47 y3 0 x47 0 0.425270206763784
Gyc3_48 y3 0 x48 0 0.419348401511974
Gyc3_49 y3 0 x49 0 0.330437217828842
Gyc3_50 y3 0 x50 0 0.434108023208343
Gyc3_51 y3 0 x51 0 0.380738404304794
Gyc3_52 y3 0 x52 0 0.313790022685357
Gyc3_53 y3 0 x53 0 -0.469306333361722
Gyc3_54 y3 0 x54 0 -0.625738619601835
Gyc3_55 y3 0 x55 0 1
Gyc3_56 y3 0 x56 0 1
Gyc3_57 y3 0 x57 0 -1
Gyc3_58 y3 0 x58 0 -1
Gyc3_59 y3 0 x59 0 1
Gyc3_60 y3 0 x60 0 0.566884191602458
Gyc3_61 y3 0 x61 0 1
Gyc3_62 y3 0 x62 0 -1
Gyc3_63 y3 0 x63 0 0.782942634623537
Gyc3_64 y3 0 x64 0 0.179559279189002
Gyc3_65 y3 0 x65 0 -0.0992057245022242
Gyc3_66 y3 0 x66 0 0.641384090293352
Gyc3_67 y3 0 x67 0 -1
Gyc3_68 y3 0 x68 0 -1
Gyc3_69 y3 0 x69 0 -0.018776795674913
Gyc3_70 y3 0 x70 0 0.0328238371067473
Gyc3_71 y3 0 x71 0 1
Gyc3_72 y3 0 x72 0 1
Gyc3_73 y3 0 x73 0 -1
Gyc3_74 y3 0 x74 0 0.306387753106672
Gyc3_75 y3 0 x75 0 -0.115618212400027
Gyc3_76 y3 0 x76 0 -0.525425155381433
Gyc3_77 y3 0 x77 0 -1
Gyc3_78 y3 0 x78 0 1
Gyc3_79 y3 0 x79 0 0.191374066155789
Gyc3_80 y3 0 x80 0 0.63058503678395
Gyc3_81 y3 0 x81 0 -0.295387547309993
.ENDS
