* Equivalent circuit model for E:\touchstone_files\15p.ckt
.SUBCKT 15p po1 po2
Vsp1 po1 p1 0
Vsr1 p1 pr1 0
Rp1 pr1 0 50
Ru1 u1 0 50
Fr1 u1 0 Vsr1 -1
Fu1 u1 0 Vsp1 -1
Ry1 y1 0 1
Gy1 p1 0 y1 0 -0.02
Vsp2 po2 p2 0
Vsr2 p2 pr2 0
Rp2 pr2 0 50
Ru2 u2 0 50
Fr2 u2 0 Vsr2 -1
Fu2 u2 0 Vsp2 -1
Ry2 y2 0 1
Gy2 p2 0 y2 0 -0.02
Rx1 x1 0 1
Fxc1_2 x1 0 Vx2 0.150262594888616
Cx1 x1 xm1 1.51671056394881e-13
Vx1 xm1 0 0
Gx1_1 x1 0 u1 0 -0.115687630135364
Rx2 x2 0 1
Fxc2_1 x2 0 Vx1 -7.58798837718887
Cx2 x2 xm2 1.51671056394881e-13
Vx2 xm2 0 0
Gx2_1 x2 0 u1 0 0.87783639285167
Rx3 x3 0 1
Cx3 x3 0 5.83463769623474e-12
Gx3_1 x3 0 u1 0 -0.0103777039075621
Rx4 x4 0 1
Fxc4_5 x4 0 Vx5 0.150265066712227
Cx4 x4 xm4 1.51671056394881e-13
Vx4 xm4 0 0
Gx4_2 x4 0 u2 0 -0.115688609541307
Rx5 x5 0 1
Fxc5_4 x5 0 Vx4 -7.58786355663518
Cx5 x5 xm5 1.51671056394881e-13
Vx5 xm5 0 0
Gx5_2 x5 0 u2 0 0.877829384256278
Rx6 x6 0 1
Cx6 x6 0 5.83463769623474e-12
Gx6_2 x6 0 u2 0 -0.0103831778540376
Gyc1_1 y1 0 x1 0 0.433699392530763
Gyc1_2 y1 0 x2 0 0.059710285114995
Gyc1_3 y1 0 x3 0 0.100139437847313
Gyc1_4 y1 0 x4 0 -1
Gyc1_5 y1 0 x5 0 1
Gyc1_6 y1 0 x6 0 -1
Gyc2_1 y2 0 x1 0 -1
Gyc2_2 y2 0 x2 0 1
Gyc2_3 y2 0 x3 0 -1
Gyc2_4 y2 0 x4 0 0.431614456801147
Gyc2_5 y2 0 x5 0 0.0594703747896991
Gyc2_6 y2 0 x6 0 0.102894430086451
.ENDS
