* Equivalent circuit model for E:\touchstone_files\35p.ckt
.SUBCKT 35p po1 po2
Vsp1 po1 p1 0
Vsr1 p1 pr1 0
Rp1 pr1 0 50
Ru1 u1 0 50
Fr1 u1 0 Vsr1 -1
Fu1 u1 0 Vsp1 -1
Ry1 y1 0 1
Gy1 p1 0 y1 0 -0.02
Vsp2 po2 p2 0
Vsr2 p2 pr2 0
Rp2 pr2 0 50
Ru2 u2 0 50
Fr2 u2 0 Vsr2 -1
Fu2 u2 0 Vsp2 -1
Ry2 y2 0 1
Gy2 p2 0 y2 0 -0.02
Rx1 x1 0 1
Fxc1_2 x1 0 Vx2 0.026745847124408
Cx1 x1 xm1 3.37735547881525e-13
Vx1 xm1 0 0
Gx1_1 x1 0 u1 0 -0.0321064425216062
Rx2 x2 0 1
Fxc2_1 x2 0 Vx1 -19.5402230749782
Cx2 x2 xm2 3.37735547881525e-13
Vx2 xm2 0 0
Gx2_1 x2 0 u1 0 0.62736704901615
Rx3 x3 0 1
Fxc3_4 x3 0 Vx4 1.61526802726054
Cx3 x3 xm3 1.20016649303951e-13
Vx3 xm3 0 0
Gx3_1 x3 0 u1 0 -0.164975846668597
Rx4 x4 0 1
Fxc4_3 x4 0 Vx3 -3.17244719353881
Cx4 x4 xm4 1.20016649303951e-13
Vx4 xm4 0 0
Gx4_1 x4 0 u1 0 0.523377161765479
Rx5 x5 0 1
Cx5 x5 0 6.21233205378623e-12
Gx5_1 x5 0 u1 0 -0.00684540393607525
Rx6 x6 0 1
Fxc6_7 x6 0 Vx7 0.0251149973201163
Cx6 x6 xm6 3.37735547881525e-13
Vx6 xm6 0 0
Gx6_2 x6 0 u2 0 -0.0301483637269103
Rx7 x7 0 1
Fxc7_6 x7 0 Vx6 -20.8090732592512
Cx7 x7 xm7 3.37735547881525e-13
Vx7 xm7 0 0
Gx7_2 x7 0 u2 0 0.627359509439828
Rx8 x8 0 1
Fxc8_9 x8 0 Vx9 1.61506222033934
Cx8 x8 xm8 1.20016649303951e-13
Vx8 xm8 0 0
Gx8_2 x8 0 u2 0 -0.164972337931783
Rx9 x9 0 1
Fxc9_8 x9 0 Vx8 -3.17285145758595
Cx9 x9 xm9 1.20016649303951e-13
Vx9 xm9 0 0
Gx9_2 x9 0 u2 0 0.523432722868219
Rx10 x10 0 1
Cx10 x10 0 6.21233205378623e-12
Gx10_2 x10 0 u2 0 -0.00685463725318149
Gyc1_1 y1 0 x1 0 1
Gyc1_2 y1 0 x2 0 0.0791315224088337
Gyc1_3 y1 0 x3 0 -0.0257838220418004
Gyc1_4 y1 0 x4 0 -0.0305150867921971
Gyc1_5 y1 0 x5 0 0.455015138591104
Gyc1_6 y1 0 x6 0 -0.179521917823964
Gyc1_7 y1 0 x7 0 1
Gyc1_8 y1 0 x8 0 1
Gyc1_9 y1 0 x9 0 1
Gyc1_10 y1 0 x10 0 -1
Gyc2_1 y2 0 x1 0 -0.170528070609993
Gyc2_2 y2 0 x2 0 1
Gyc2_3 y2 0 x3 0 1
Gyc2_4 y2 0 x4 0 1
Gyc2_5 y2 0 x5 0 -1
Gyc2_6 y2 0 x6 0 1
Gyc2_7 y2 0 x7 0 0.0784075317911112
Gyc2_8 y2 0 x8 0 -0.0257481080632151
Gyc2_9 y2 0 x9 0 -0.0334501505266849
Gyc2_10 y2 0 x10 0 0.449603020084359
.ENDS
